`ifndef __CORE__
`define __CORE__

`include "VGASyncGen.vh"

`endif
